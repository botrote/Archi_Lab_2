module alu (
	input [`WORD_SIZE-1:0] address,
	input [`WORD_SIZE-1:0] write_data,

	input signal_MemToRead,
	input signal_MemWrite,
	input clk

	output [`WORD_SIZE-1:0] read_data
);

	assign read_data = 

	integer i;
	always @ (posedge clk or posedge reset_n) begin
		if(reset_n)
			for(i = 0; i < ; i = i + 1)

		else


endmodule

//NOT REQUIRED